-- Sumador completo de un bit
-- Recibe 3 bits: a, b y el acarreo de entrada cin
-- Retorna el bit de sumatoria (sum) y el acarreo de salida cout
LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity BIT_ADDER_1 is
	port( a, b, cin         : in  STD_LOGIC;
	      sum, cout         : out STD_LOGIC );
end BIT_ADDER_1;

architecture BHV of BIT_ADDER_1 is
begin
	
	-- Calculate the sum of the 1-BIT adder.
	sum <=  (a xor b) xor cin;
	-- Calculates the carry out of the 1-BIT adder.
	cout <= (a and b) or (cin and (a xor b));
end BHV;





-- Sumador completo de 4 bits
-- Utiliza sumadores de 1 bit interconectando sus salidas y acarreos con nuevas entradas
-- Recibe dos vectores de 4 bits a y b. Además recibe el acarreo de entrada
-- Retorna 4 bits de sumatoria (sum) y el acarreo de salida cout

LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity adder4_aux is
	port( a, b		: in	STD_LOGIC_VECTOR(3 downto 0);
			cin      : in STD_LOGIC;
	      ans		: out	STD_LOGIC_VECTOR(3 downto 0);
	      cout		: out	STD_LOGIC);
end adder4_aux;



architecture STRUCTURE of adder4_aux is


component BIT_ADDER_1
	port( a, b, cin		: in  STD_LOGIC;
	      sum, cout		: out STD_LOGIC );
end component;



-- Utilización de cada sumador de 1 bit por medio de señales que pasan la información
signal c1, c2, c3 : STD_LOGIC;
begin

b_adder0: BIT_ADDER_1 port map (a(0), b(0), cin, ans(0), c1);
b_adder1: BIT_ADDER_1 port map (a(1), b(1), c1, ans(1), c2);
b_adder2: BIT_ADDER_1 port map (a(2), b(2), c2, ans(2), c3);
b_adder3: BIT_ADDER_1 port map (a(3), b(3), c3, ans(3), cout);


END STRUCTURE;


-- Salida del módulo de 4 bits hacia dos displays
-- Utiliza un decodificador de 4 bits a 7 para ser utilizados por el display de la FPGA
LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity adder4 is
	port( a, b		: in	STD_LOGIC_VECTOR(3 downto 0);
			cin      : in STD_LOGIC;
			ans		: out	STD_LOGIC_VECTOR(3 downto 0);
			cout		: out STD_LOGIC;
	      display 	: out STD_LOGIC_VECTOR(6 downto 0);
			display_aux :out STD_LOGIC_VECTOR(6 downto 0));
end adder4;


architecture BHV of adder4 is
component adder4_aux
	port( a, b		: in	STD_LOGIC_VECTOR(3 downto 0);
			cin      : in STD_LOGIC;
	      ans		: out	STD_LOGIC_VECTOR(3 downto 0);
	      cout		: out	STD_LOGIC);
end component;

signal ans_aux, ans_aux_2  : STD_LOGIC_VECTOR(3 downto 0);
signal cout_aux : STD_LOGIC;

begin

	adder4_1 : adder4_aux port map (a, b, cin, ans_aux_2, cout_aux);
	process(ans_aux_2)
	begin
		case ans_aux_2 is
			when "0000" => display <= "1000000"; -- "0"    0000001 
			when "0001" => display <= "1111001"; -- "1"    1001111
			when "0010" => display <= "0100100"; -- "2"    0010010
			when "0011" => display <= "0110000"; -- "3" 	  0000110
			when "0100" => display <= "0011001"; -- "4"    1001100
			when "0101" => display <= "0010010"; -- "5"    0100100
			when "0110" => display <= "0000010"; -- "6"    0100000
			when "0111" => display <= "1111000"; -- "7"    0001111
			when "1000" => display <= "0000000"; -- "8"     
			when "1001" => display <= "0010000"; -- "9"    0000100
			when "1010" => display <= "0100000"; -- a      0000010
			when "1011" => display <= "0000011"; -- b
			when "1100" => display <= "1000110"; -- C      0110001
			when "1101" => display <= "0100001"; -- d      1000010
			when "1110" => display <= "0000110"; -- E
			when "1111" => display <= "0001110"; -- F
			when others => display <= "1000000"; -- "0"    0000001 
		end case;
	end process;
	
	process(cout_aux)
	begin
		case cout_aux is
			when '0' => display_aux <= "1000000"; -- "0"     
			when '1' => display_aux <= "1111001"; -- "1" 
			when others => display_aux <= "1000000"; -- "0" 
		end case;
	end process;
	ans <= ans_aux_2;
	cout <= cout_aux;
	
	
end BHV;
