module ecualizador_histograma_tb;


endmodule