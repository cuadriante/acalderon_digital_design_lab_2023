module f5(input I0, I1, I2, I3, output S4);

	assign S4 = (I3);
	
endmodule

